module bench_spi_recv_pu ();

    
endmodule